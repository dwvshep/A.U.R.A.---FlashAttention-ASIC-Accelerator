//This module computes the exponential multiplication of a scalar with a vector combinationally

module expmul_comb(
    //Data signals
    input INT_T a_in,
    input INT_T b_in,
    input STAR_VECTOR_T v_in,
    output STAR_VECTOR_T v_out
);

    //output is combinational
    always_comb begin

    end

endmodule