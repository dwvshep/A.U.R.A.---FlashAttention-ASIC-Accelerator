module dot_product(
    //Handshake signals
    input vld_in,
    input rdy_in,
    output vld_out,
    output rdy_out,

    //Data signals
    input Q_VECTOR_T q_in,
    input K_VECTOR_T k_in,
);


endmodule