module memory_controller(
    input clk,
    input rst,

    input logic Q_sram_ready,
    output logic ctrl_ready,
    
);


endmodule