module controller(

);


endmodule