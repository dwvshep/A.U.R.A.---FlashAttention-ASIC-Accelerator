module memory_controller(

);


endmodule